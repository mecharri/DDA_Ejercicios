always@(posedge clock) begin
  coeff[0]  <= 8'd0;
  coeff[1]  <= 8'd0;
  coeff[2]  <= 8'd1;
  coeff[3]  <= 8'd4;
  coeff[4]  <= 8'd10;
  coeff[5]  <= 8'd16;
  coeff[6]  <= 8'd21;
  coeff[7]  <= 8'd24;
  coeff[8]  <= 8'd21;
  coeff[9]  <= 8'd16;
  coeff[10]  <= 8'd10;
  coeff[11]  <= 8'd4;
  coeff[12]  <= 8'd1;
  coeff[13]  <= 8'd0;
  coeff[14]  <= 8'd0;
end